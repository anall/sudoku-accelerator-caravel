magic
tech sky130A
magscale 1 2
timestamp 1634053839
<< obsli1 >>
rect 1104 1377 165968 167025
<< obsm1 >>
rect 106 824 166598 167056
<< metal2 >>
rect 662 168478 718 169278
rect 2042 168478 2098 169278
rect 3514 168478 3570 169278
rect 4894 168478 4950 169278
rect 6366 168478 6422 169278
rect 7838 168478 7894 169278
rect 9218 168478 9274 169278
rect 10690 168478 10746 169278
rect 12162 168478 12218 169278
rect 13542 168478 13598 169278
rect 15014 168478 15070 169278
rect 16486 168478 16542 169278
rect 17866 168478 17922 169278
rect 19338 168478 19394 169278
rect 20810 168478 20866 169278
rect 22190 168478 22246 169278
rect 23662 168478 23718 169278
rect 25134 168478 25190 169278
rect 26514 168478 26570 169278
rect 27986 168478 28042 169278
rect 29458 168478 29514 169278
rect 30838 168478 30894 169278
rect 32310 168478 32366 169278
rect 33782 168478 33838 169278
rect 35162 168478 35218 169278
rect 36634 168478 36690 169278
rect 38106 168478 38162 169278
rect 39486 168478 39542 169278
rect 40958 168478 41014 169278
rect 42430 168478 42486 169278
rect 43810 168478 43866 169278
rect 45282 168478 45338 169278
rect 46754 168478 46810 169278
rect 48134 168478 48190 169278
rect 49606 168478 49662 169278
rect 51078 168478 51134 169278
rect 52458 168478 52514 169278
rect 53930 168478 53986 169278
rect 55402 168478 55458 169278
rect 56782 168478 56838 169278
rect 58254 168478 58310 169278
rect 59726 168478 59782 169278
rect 61106 168478 61162 169278
rect 62578 168478 62634 169278
rect 64050 168478 64106 169278
rect 65430 168478 65486 169278
rect 66902 168478 66958 169278
rect 68374 168478 68430 169278
rect 69754 168478 69810 169278
rect 71226 168478 71282 169278
rect 72698 168478 72754 169278
rect 74078 168478 74134 169278
rect 75550 168478 75606 169278
rect 77022 168478 77078 169278
rect 78402 168478 78458 169278
rect 79874 168478 79930 169278
rect 81346 168478 81402 169278
rect 82726 168478 82782 169278
rect 84198 168478 84254 169278
rect 85670 168478 85726 169278
rect 87050 168478 87106 169278
rect 88522 168478 88578 169278
rect 89994 168478 90050 169278
rect 91374 168478 91430 169278
rect 92846 168478 92902 169278
rect 94318 168478 94374 169278
rect 95698 168478 95754 169278
rect 97170 168478 97226 169278
rect 98642 168478 98698 169278
rect 100022 168478 100078 169278
rect 101494 168478 101550 169278
rect 102966 168478 103022 169278
rect 104346 168478 104402 169278
rect 105818 168478 105874 169278
rect 107290 168478 107346 169278
rect 108670 168478 108726 169278
rect 110142 168478 110198 169278
rect 111614 168478 111670 169278
rect 112994 168478 113050 169278
rect 114466 168478 114522 169278
rect 115938 168478 115994 169278
rect 117318 168478 117374 169278
rect 118790 168478 118846 169278
rect 120262 168478 120318 169278
rect 121642 168478 121698 169278
rect 123114 168478 123170 169278
rect 124586 168478 124642 169278
rect 125966 168478 126022 169278
rect 127438 168478 127494 169278
rect 128910 168478 128966 169278
rect 130290 168478 130346 169278
rect 131762 168478 131818 169278
rect 133234 168478 133290 169278
rect 134614 168478 134670 169278
rect 136086 168478 136142 169278
rect 137558 168478 137614 169278
rect 138938 168478 138994 169278
rect 140410 168478 140466 169278
rect 141882 168478 141938 169278
rect 143262 168478 143318 169278
rect 144734 168478 144790 169278
rect 146206 168478 146262 169278
rect 147586 168478 147642 169278
rect 149058 168478 149114 169278
rect 150530 168478 150586 169278
rect 151910 168478 151966 169278
rect 153382 168478 153438 169278
rect 154854 168478 154910 169278
rect 156234 168478 156290 169278
rect 157706 168478 157762 169278
rect 159178 168478 159234 169278
rect 160558 168478 160614 169278
rect 162030 168478 162086 169278
rect 163502 168478 163558 169278
rect 164882 168478 164938 169278
rect 166354 168478 166410 169278
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61474 0 61530 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89442 0 89498 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91466 0 91522 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119434 0 119490 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123206 0 123262 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155590 0 155646 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159362 0 159418 800
rect 159730 0 159786 800
rect 160098 0 160154 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161110 0 161166 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162766 0 162822 800
rect 163134 0 163190 800
rect 163502 0 163558 800
rect 163778 0 163834 800
rect 164146 0 164202 800
rect 164514 0 164570 800
rect 164882 0 164938 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
<< obsm2 >>
rect 18 168422 606 168586
rect 774 168422 1986 168586
rect 2154 168422 3458 168586
rect 3626 168422 4838 168586
rect 5006 168422 6310 168586
rect 6478 168422 7782 168586
rect 7950 168422 9162 168586
rect 9330 168422 10634 168586
rect 10802 168422 12106 168586
rect 12274 168422 13486 168586
rect 13654 168422 14958 168586
rect 15126 168422 16430 168586
rect 16598 168422 17810 168586
rect 17978 168422 19282 168586
rect 19450 168422 20754 168586
rect 20922 168422 22134 168586
rect 22302 168422 23606 168586
rect 23774 168422 25078 168586
rect 25246 168422 26458 168586
rect 26626 168422 27930 168586
rect 28098 168422 29402 168586
rect 29570 168422 30782 168586
rect 30950 168422 32254 168586
rect 32422 168422 33726 168586
rect 33894 168422 35106 168586
rect 35274 168422 36578 168586
rect 36746 168422 38050 168586
rect 38218 168422 39430 168586
rect 39598 168422 40902 168586
rect 41070 168422 42374 168586
rect 42542 168422 43754 168586
rect 43922 168422 45226 168586
rect 45394 168422 46698 168586
rect 46866 168422 48078 168586
rect 48246 168422 49550 168586
rect 49718 168422 51022 168586
rect 51190 168422 52402 168586
rect 52570 168422 53874 168586
rect 54042 168422 55346 168586
rect 55514 168422 56726 168586
rect 56894 168422 58198 168586
rect 58366 168422 59670 168586
rect 59838 168422 61050 168586
rect 61218 168422 62522 168586
rect 62690 168422 63994 168586
rect 64162 168422 65374 168586
rect 65542 168422 66846 168586
rect 67014 168422 68318 168586
rect 68486 168422 69698 168586
rect 69866 168422 71170 168586
rect 71338 168422 72642 168586
rect 72810 168422 74022 168586
rect 74190 168422 75494 168586
rect 75662 168422 76966 168586
rect 77134 168422 78346 168586
rect 78514 168422 79818 168586
rect 79986 168422 81290 168586
rect 81458 168422 82670 168586
rect 82838 168422 84142 168586
rect 84310 168422 85614 168586
rect 85782 168422 86994 168586
rect 87162 168422 88466 168586
rect 88634 168422 89938 168586
rect 90106 168422 91318 168586
rect 91486 168422 92790 168586
rect 92958 168422 94262 168586
rect 94430 168422 95642 168586
rect 95810 168422 97114 168586
rect 97282 168422 98586 168586
rect 98754 168422 99966 168586
rect 100134 168422 101438 168586
rect 101606 168422 102910 168586
rect 103078 168422 104290 168586
rect 104458 168422 105762 168586
rect 105930 168422 107234 168586
rect 107402 168422 108614 168586
rect 108782 168422 110086 168586
rect 110254 168422 111558 168586
rect 111726 168422 112938 168586
rect 113106 168422 114410 168586
rect 114578 168422 115882 168586
rect 116050 168422 117262 168586
rect 117430 168422 118734 168586
rect 118902 168422 120206 168586
rect 120374 168422 121586 168586
rect 121754 168422 123058 168586
rect 123226 168422 124530 168586
rect 124698 168422 125910 168586
rect 126078 168422 127382 168586
rect 127550 168422 128854 168586
rect 129022 168422 130234 168586
rect 130402 168422 131706 168586
rect 131874 168422 133178 168586
rect 133346 168422 134558 168586
rect 134726 168422 136030 168586
rect 136198 168422 137502 168586
rect 137670 168422 138882 168586
rect 139050 168422 140354 168586
rect 140522 168422 141826 168586
rect 141994 168422 143206 168586
rect 143374 168422 144678 168586
rect 144846 168422 146150 168586
rect 146318 168422 147530 168586
rect 147698 168422 149002 168586
rect 149170 168422 150474 168586
rect 150642 168422 151854 168586
rect 152022 168422 153326 168586
rect 153494 168422 154798 168586
rect 154966 168422 156178 168586
rect 156346 168422 157650 168586
rect 157818 168422 159122 168586
rect 159290 168422 160502 168586
rect 160670 168422 161974 168586
rect 162142 168422 163446 168586
rect 163614 168422 164826 168586
rect 164994 168422 166298 168586
rect 166466 168422 166592 168586
rect 18 856 166592 168422
rect 18 734 54 856
rect 222 734 330 856
rect 498 734 698 856
rect 866 734 1066 856
rect 1234 734 1342 856
rect 1510 734 1710 856
rect 1878 734 2078 856
rect 2246 734 2354 856
rect 2522 734 2722 856
rect 2890 734 3090 856
rect 3258 734 3458 856
rect 3626 734 3734 856
rect 3902 734 4102 856
rect 4270 734 4470 856
rect 4638 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6126 856
rect 6294 734 6494 856
rect 6662 734 6862 856
rect 7030 734 7138 856
rect 7306 734 7506 856
rect 7674 734 7874 856
rect 8042 734 8150 856
rect 8318 734 8518 856
rect 8686 734 8886 856
rect 9054 734 9254 856
rect 9422 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10266 856
rect 10434 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 11922 856
rect 12090 734 12290 856
rect 12458 734 12658 856
rect 12826 734 12934 856
rect 13102 734 13302 856
rect 13470 734 13670 856
rect 13838 734 14038 856
rect 14206 734 14314 856
rect 14482 734 14682 856
rect 14850 734 15050 856
rect 15218 734 15326 856
rect 15494 734 15694 856
rect 15862 734 16062 856
rect 16230 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17718 856
rect 17886 734 18086 856
rect 18254 734 18454 856
rect 18622 734 18730 856
rect 18898 734 19098 856
rect 19266 734 19466 856
rect 19634 734 19834 856
rect 20002 734 20110 856
rect 20278 734 20478 856
rect 20646 734 20846 856
rect 21014 734 21122 856
rect 21290 734 21490 856
rect 21658 734 21858 856
rect 22026 734 22226 856
rect 22394 734 22502 856
rect 22670 734 22870 856
rect 23038 734 23238 856
rect 23406 734 23514 856
rect 23682 734 23882 856
rect 24050 734 24250 856
rect 24418 734 24526 856
rect 24694 734 24894 856
rect 25062 734 25262 856
rect 25430 734 25630 856
rect 25798 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27654 856
rect 27822 734 28022 856
rect 28190 734 28298 856
rect 28466 734 28666 856
rect 28834 734 29034 856
rect 29202 734 29310 856
rect 29478 734 29678 856
rect 29846 734 30046 856
rect 30214 734 30414 856
rect 30582 734 30690 856
rect 30858 734 31058 856
rect 31226 734 31426 856
rect 31594 734 31702 856
rect 31870 734 32070 856
rect 32238 734 32438 856
rect 32606 734 32714 856
rect 32882 734 33082 856
rect 33250 734 33450 856
rect 33618 734 33818 856
rect 33986 734 34094 856
rect 34262 734 34462 856
rect 34630 734 34830 856
rect 34998 734 35106 856
rect 35274 734 35474 856
rect 35642 734 35842 856
rect 36010 734 36210 856
rect 36378 734 36486 856
rect 36654 734 36854 856
rect 37022 734 37222 856
rect 37390 734 37498 856
rect 37666 734 37866 856
rect 38034 734 38234 856
rect 38402 734 38602 856
rect 38770 734 38878 856
rect 39046 734 39246 856
rect 39414 734 39614 856
rect 39782 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40626 856
rect 40794 734 40902 856
rect 41070 734 41270 856
rect 41438 734 41638 856
rect 41806 734 42006 856
rect 42174 734 42282 856
rect 42450 734 42650 856
rect 42818 734 43018 856
rect 43186 734 43294 856
rect 43462 734 43662 856
rect 43830 734 44030 856
rect 44198 734 44398 856
rect 44566 734 44674 856
rect 44842 734 45042 856
rect 45210 734 45410 856
rect 45578 734 45686 856
rect 45854 734 46054 856
rect 46222 734 46422 856
rect 46590 734 46790 856
rect 46958 734 47066 856
rect 47234 734 47434 856
rect 47602 734 47802 856
rect 47970 734 48078 856
rect 48246 734 48446 856
rect 48614 734 48814 856
rect 48982 734 49090 856
rect 49258 734 49458 856
rect 49626 734 49826 856
rect 49994 734 50194 856
rect 50362 734 50470 856
rect 50638 734 50838 856
rect 51006 734 51206 856
rect 51374 734 51482 856
rect 51650 734 51850 856
rect 52018 734 52218 856
rect 52386 734 52586 856
rect 52754 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53874 856
rect 54042 734 54242 856
rect 54410 734 54610 856
rect 54778 734 54978 856
rect 55146 734 55254 856
rect 55422 734 55622 856
rect 55790 734 55990 856
rect 56158 734 56266 856
rect 56434 734 56634 856
rect 56802 734 57002 856
rect 57170 734 57278 856
rect 57446 734 57646 856
rect 57814 734 58014 856
rect 58182 734 58382 856
rect 58550 734 58658 856
rect 58826 734 59026 856
rect 59194 734 59394 856
rect 59562 734 59670 856
rect 59838 734 60038 856
rect 60206 734 60406 856
rect 60574 734 60774 856
rect 60942 734 61050 856
rect 61218 734 61418 856
rect 61586 734 61786 856
rect 61954 734 62062 856
rect 62230 734 62430 856
rect 62598 734 62798 856
rect 62966 734 63166 856
rect 63334 734 63442 856
rect 63610 734 63810 856
rect 63978 734 64178 856
rect 64346 734 64454 856
rect 64622 734 64822 856
rect 64990 734 65190 856
rect 65358 734 65466 856
rect 65634 734 65834 856
rect 66002 734 66202 856
rect 66370 734 66570 856
rect 66738 734 66846 856
rect 67014 734 67214 856
rect 67382 734 67582 856
rect 67750 734 67858 856
rect 68026 734 68226 856
rect 68394 734 68594 856
rect 68762 734 68962 856
rect 69130 734 69238 856
rect 69406 734 69606 856
rect 69774 734 69974 856
rect 70142 734 70250 856
rect 70418 734 70618 856
rect 70786 734 70986 856
rect 71154 734 71354 856
rect 71522 734 71630 856
rect 71798 734 71998 856
rect 72166 734 72366 856
rect 72534 734 72642 856
rect 72810 734 73010 856
rect 73178 734 73378 856
rect 73546 734 73654 856
rect 73822 734 74022 856
rect 74190 734 74390 856
rect 74558 734 74758 856
rect 74926 734 75034 856
rect 75202 734 75402 856
rect 75570 734 75770 856
rect 75938 734 76046 856
rect 76214 734 76414 856
rect 76582 734 76782 856
rect 76950 734 77150 856
rect 77318 734 77426 856
rect 77594 734 77794 856
rect 77962 734 78162 856
rect 78330 734 78438 856
rect 78606 734 78806 856
rect 78974 734 79174 856
rect 79342 734 79542 856
rect 79710 734 79818 856
rect 79986 734 80186 856
rect 80354 734 80554 856
rect 80722 734 80830 856
rect 80998 734 81198 856
rect 81366 734 81566 856
rect 81734 734 81842 856
rect 82010 734 82210 856
rect 82378 734 82578 856
rect 82746 734 82946 856
rect 83114 734 83222 856
rect 83390 734 83590 856
rect 83758 734 83958 856
rect 84126 734 84234 856
rect 84402 734 84602 856
rect 84770 734 84970 856
rect 85138 734 85338 856
rect 85506 734 85614 856
rect 85782 734 85982 856
rect 86150 734 86350 856
rect 86518 734 86626 856
rect 86794 734 86994 856
rect 87162 734 87362 856
rect 87530 734 87638 856
rect 87806 734 88006 856
rect 88174 734 88374 856
rect 88542 734 88742 856
rect 88910 734 89018 856
rect 89186 734 89386 856
rect 89554 734 89754 856
rect 89922 734 90030 856
rect 90198 734 90398 856
rect 90566 734 90766 856
rect 90934 734 91134 856
rect 91302 734 91410 856
rect 91578 734 91778 856
rect 91946 734 92146 856
rect 92314 734 92422 856
rect 92590 734 92790 856
rect 92958 734 93158 856
rect 93326 734 93526 856
rect 93694 734 93802 856
rect 93970 734 94170 856
rect 94338 734 94538 856
rect 94706 734 94814 856
rect 94982 734 95182 856
rect 95350 734 95550 856
rect 95718 734 95826 856
rect 95994 734 96194 856
rect 96362 734 96562 856
rect 96730 734 96930 856
rect 97098 734 97206 856
rect 97374 734 97574 856
rect 97742 734 97942 856
rect 98110 734 98218 856
rect 98386 734 98586 856
rect 98754 734 98954 856
rect 99122 734 99322 856
rect 99490 734 99598 856
rect 99766 734 99966 856
rect 100134 734 100334 856
rect 100502 734 100610 856
rect 100778 734 100978 856
rect 101146 734 101346 856
rect 101514 734 101714 856
rect 101882 734 101990 856
rect 102158 734 102358 856
rect 102526 734 102726 856
rect 102894 734 103002 856
rect 103170 734 103370 856
rect 103538 734 103738 856
rect 103906 734 104014 856
rect 104182 734 104382 856
rect 104550 734 104750 856
rect 104918 734 105118 856
rect 105286 734 105394 856
rect 105562 734 105762 856
rect 105930 734 106130 856
rect 106298 734 106406 856
rect 106574 734 106774 856
rect 106942 734 107142 856
rect 107310 734 107510 856
rect 107678 734 107786 856
rect 107954 734 108154 856
rect 108322 734 108522 856
rect 108690 734 108798 856
rect 108966 734 109166 856
rect 109334 734 109534 856
rect 109702 734 109902 856
rect 110070 734 110178 856
rect 110346 734 110546 856
rect 110714 734 110914 856
rect 111082 734 111190 856
rect 111358 734 111558 856
rect 111726 734 111926 856
rect 112094 734 112202 856
rect 112370 734 112570 856
rect 112738 734 112938 856
rect 113106 734 113306 856
rect 113474 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114318 856
rect 114486 734 114594 856
rect 114762 734 114962 856
rect 115130 734 115330 856
rect 115498 734 115698 856
rect 115866 734 115974 856
rect 116142 734 116342 856
rect 116510 734 116710 856
rect 116878 734 116986 856
rect 117154 734 117354 856
rect 117522 734 117722 856
rect 117890 734 118090 856
rect 118258 734 118366 856
rect 118534 734 118734 856
rect 118902 734 119102 856
rect 119270 734 119378 856
rect 119546 734 119746 856
rect 119914 734 120114 856
rect 120282 734 120390 856
rect 120558 734 120758 856
rect 120926 734 121126 856
rect 121294 734 121494 856
rect 121662 734 121770 856
rect 121938 734 122138 856
rect 122306 734 122506 856
rect 122674 734 122782 856
rect 122950 734 123150 856
rect 123318 734 123518 856
rect 123686 734 123886 856
rect 124054 734 124162 856
rect 124330 734 124530 856
rect 124698 734 124898 856
rect 125066 734 125174 856
rect 125342 734 125542 856
rect 125710 734 125910 856
rect 126078 734 126278 856
rect 126446 734 126554 856
rect 126722 734 126922 856
rect 127090 734 127290 856
rect 127458 734 127566 856
rect 127734 734 127934 856
rect 128102 734 128302 856
rect 128470 734 128578 856
rect 128746 734 128946 856
rect 129114 734 129314 856
rect 129482 734 129682 856
rect 129850 734 129958 856
rect 130126 734 130326 856
rect 130494 734 130694 856
rect 130862 734 130970 856
rect 131138 734 131338 856
rect 131506 734 131706 856
rect 131874 734 132074 856
rect 132242 734 132350 856
rect 132518 734 132718 856
rect 132886 734 133086 856
rect 133254 734 133362 856
rect 133530 734 133730 856
rect 133898 734 134098 856
rect 134266 734 134466 856
rect 134634 734 134742 856
rect 134910 734 135110 856
rect 135278 734 135478 856
rect 135646 734 135754 856
rect 135922 734 136122 856
rect 136290 734 136490 856
rect 136658 734 136766 856
rect 136934 734 137134 856
rect 137302 734 137502 856
rect 137670 734 137870 856
rect 138038 734 138146 856
rect 138314 734 138514 856
rect 138682 734 138882 856
rect 139050 734 139158 856
rect 139326 734 139526 856
rect 139694 734 139894 856
rect 140062 734 140262 856
rect 140430 734 140538 856
rect 140706 734 140906 856
rect 141074 734 141274 856
rect 141442 734 141550 856
rect 141718 734 141918 856
rect 142086 734 142286 856
rect 142454 734 142654 856
rect 142822 734 142930 856
rect 143098 734 143298 856
rect 143466 734 143666 856
rect 143834 734 143942 856
rect 144110 734 144310 856
rect 144478 734 144678 856
rect 144846 734 144954 856
rect 145122 734 145322 856
rect 145490 734 145690 856
rect 145858 734 146058 856
rect 146226 734 146334 856
rect 146502 734 146702 856
rect 146870 734 147070 856
rect 147238 734 147346 856
rect 147514 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148450 856
rect 148618 734 148726 856
rect 148894 734 149094 856
rect 149262 734 149462 856
rect 149630 734 149738 856
rect 149906 734 150106 856
rect 150274 734 150474 856
rect 150642 734 150842 856
rect 151010 734 151118 856
rect 151286 734 151486 856
rect 151654 734 151854 856
rect 152022 734 152130 856
rect 152298 734 152498 856
rect 152666 734 152866 856
rect 153034 734 153142 856
rect 153310 734 153510 856
rect 153678 734 153878 856
rect 154046 734 154246 856
rect 154414 734 154522 856
rect 154690 734 154890 856
rect 155058 734 155258 856
rect 155426 734 155534 856
rect 155702 734 155902 856
rect 156070 734 156270 856
rect 156438 734 156638 856
rect 156806 734 156914 856
rect 157082 734 157282 856
rect 157450 734 157650 856
rect 157818 734 157926 856
rect 158094 734 158294 856
rect 158462 734 158662 856
rect 158830 734 159030 856
rect 159198 734 159306 856
rect 159474 734 159674 856
rect 159842 734 160042 856
rect 160210 734 160318 856
rect 160486 734 160686 856
rect 160854 734 161054 856
rect 161222 734 161330 856
rect 161498 734 161698 856
rect 161866 734 162066 856
rect 162234 734 162434 856
rect 162602 734 162710 856
rect 162878 734 163078 856
rect 163246 734 163446 856
rect 163614 734 163722 856
rect 163890 734 164090 856
rect 164258 734 164458 856
rect 164626 734 164826 856
rect 164994 734 165102 856
rect 165270 734 165470 856
rect 165638 734 165838 856
rect 166006 734 166114 856
rect 166282 734 166482 856
<< metal3 >>
rect 166334 126896 167134 127016
rect 166334 42304 167134 42424
<< obsm3 >>
rect 13 127096 166334 167041
rect 13 126816 166254 127096
rect 13 42504 166334 126816
rect 13 42224 166254 42504
rect 13 2143 166334 42224
<< metal4 >>
rect 4208 2128 4528 167056
rect 19568 2128 19888 167056
rect 34928 2128 35248 167056
rect 50288 2128 50608 167056
rect 65648 2128 65968 167056
rect 81008 2128 81328 167056
rect 96368 2128 96688 167056
rect 111728 2128 112048 167056
rect 127088 2128 127408 167056
rect 142448 2128 142768 167056
rect 157808 2128 158128 167056
<< obsm4 >>
rect 5027 2347 19488 166565
rect 19968 2347 34848 166565
rect 35328 2347 50208 166565
rect 50688 2347 65568 166565
rect 66048 2347 80928 166565
rect 81408 2347 96288 166565
rect 96768 2347 111648 166565
rect 112128 2347 127008 166565
rect 127488 2347 142368 166565
rect 142848 2347 157728 166565
rect 158208 2347 163701 166565
<< labels >>
rlabel metal2 s 662 168478 718 169278 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43810 168478 43866 169278 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 48134 168478 48190 169278 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 52458 168478 52514 169278 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 56782 168478 56838 169278 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 61106 168478 61162 169278 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 65430 168478 65486 169278 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 69754 168478 69810 169278 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 74078 168478 74134 169278 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 78402 168478 78458 169278 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 82726 168478 82782 169278 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4894 168478 4950 169278 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 87050 168478 87106 169278 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 91374 168478 91430 169278 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 95698 168478 95754 169278 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 100022 168478 100078 169278 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 104346 168478 104402 169278 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 108670 168478 108726 169278 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 112994 168478 113050 169278 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 117318 168478 117374 169278 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 121642 168478 121698 169278 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 125966 168478 126022 169278 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9218 168478 9274 169278 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 130290 168478 130346 169278 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 134614 168478 134670 169278 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 138938 168478 138994 169278 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 143262 168478 143318 169278 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 147586 168478 147642 169278 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 151910 168478 151966 169278 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 156234 168478 156290 169278 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 160558 168478 160614 169278 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13542 168478 13598 169278 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17866 168478 17922 169278 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 22190 168478 22246 169278 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26514 168478 26570 169278 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30838 168478 30894 169278 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 35162 168478 35218 169278 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 39486 168478 39542 169278 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 168478 2098 169278 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 45282 168478 45338 169278 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 49606 168478 49662 169278 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53930 168478 53986 169278 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 58254 168478 58310 169278 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 62578 168478 62634 169278 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 66902 168478 66958 169278 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 71226 168478 71282 169278 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 75550 168478 75606 169278 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 79874 168478 79930 169278 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 84198 168478 84254 169278 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6366 168478 6422 169278 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 88522 168478 88578 169278 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 92846 168478 92902 169278 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 97170 168478 97226 169278 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 101494 168478 101550 169278 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 105818 168478 105874 169278 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 110142 168478 110198 169278 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 114466 168478 114522 169278 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 118790 168478 118846 169278 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 123114 168478 123170 169278 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 127438 168478 127494 169278 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10690 168478 10746 169278 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 131762 168478 131818 169278 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 136086 168478 136142 169278 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 140410 168478 140466 169278 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 144734 168478 144790 169278 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 149058 168478 149114 169278 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 153382 168478 153438 169278 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 157706 168478 157762 169278 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 162030 168478 162086 169278 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15014 168478 15070 169278 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19338 168478 19394 169278 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23662 168478 23718 169278 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27986 168478 28042 169278 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 32310 168478 32366 169278 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36634 168478 36690 169278 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40958 168478 41014 169278 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3514 168478 3570 169278 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46754 168478 46810 169278 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 51078 168478 51134 169278 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 55402 168478 55458 169278 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 59726 168478 59782 169278 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 64050 168478 64106 169278 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 68374 168478 68430 169278 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 72698 168478 72754 169278 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 77022 168478 77078 169278 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 81346 168478 81402 169278 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 85670 168478 85726 169278 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7838 168478 7894 169278 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 89994 168478 90050 169278 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 94318 168478 94374 169278 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 98642 168478 98698 169278 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 102966 168478 103022 169278 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 107290 168478 107346 169278 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 111614 168478 111670 169278 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 115938 168478 115994 169278 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 120262 168478 120318 169278 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 124586 168478 124642 169278 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 128910 168478 128966 169278 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12162 168478 12218 169278 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 133234 168478 133290 169278 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 137558 168478 137614 169278 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 141882 168478 141938 169278 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 146206 168478 146262 169278 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 150530 168478 150586 169278 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 154854 168478 154910 169278 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 159178 168478 159234 169278 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 163502 168478 163558 169278 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16486 168478 16542 169278 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20810 168478 20866 169278 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 25134 168478 25190 169278 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 29458 168478 29514 169278 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33782 168478 33838 169278 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 38106 168478 38162 169278 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 42430 168478 42486 169278 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_oenb[0]
port 371 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[100]
port 372 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[101]
port 373 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[102]
port 374 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[103]
port 375 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[104]
port 376 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[105]
port 377 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[106]
port 378 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[107]
port 379 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oenb[108]
port 380 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[109]
port 381 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[10]
port 382 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[110]
port 383 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_oenb[111]
port 384 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_oenb[112]
port 385 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_oenb[113]
port 386 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[114]
port 387 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[115]
port 388 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[116]
port 389 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[117]
port 390 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_oenb[118]
port 391 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[119]
port 392 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[11]
port 393 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[120]
port 394 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oenb[121]
port 395 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[122]
port 396 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[123]
port 397 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[124]
port 398 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[125]
port 399 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[126]
port 400 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_oenb[127]
port 401 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[12]
port 402 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[13]
port 403 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[14]
port 404 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[15]
port 405 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[16]
port 406 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[17]
port 407 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[18]
port 408 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[19]
port 409 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[1]
port 410 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[20]
port 411 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[21]
port 412 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[22]
port 413 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[23]
port 414 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[24]
port 415 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[25]
port 416 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[26]
port 417 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_oenb[27]
port 418 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[28]
port 419 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[29]
port 420 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[2]
port 421 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[30]
port 422 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[31]
port 423 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[32]
port 424 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[33]
port 425 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[34]
port 426 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[35]
port 427 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[36]
port 428 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[37]
port 429 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[38]
port 430 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[39]
port 431 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[3]
port 432 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[40]
port 433 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[41]
port 434 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[42]
port 435 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[43]
port 436 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[44]
port 437 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[45]
port 438 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[46]
port 439 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[47]
port 440 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[48]
port 441 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[49]
port 442 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[4]
port 443 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[50]
port 444 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[51]
port 445 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[52]
port 446 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[53]
port 447 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[54]
port 448 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[55]
port 449 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[56]
port 450 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[57]
port 451 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[58]
port 452 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[59]
port 453 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[5]
port 454 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[60]
port 455 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[61]
port 456 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[62]
port 457 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[63]
port 458 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[64]
port 459 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[65]
port 460 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[66]
port 461 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[67]
port 462 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[68]
port 463 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[69]
port 464 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[6]
port 465 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[70]
port 466 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[71]
port 467 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[72]
port 468 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[73]
port 469 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[74]
port 470 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[75]
port 471 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[76]
port 472 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oenb[77]
port 473 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[78]
port 474 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[79]
port 475 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[7]
port 476 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_oenb[80]
port 477 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[81]
port 478 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[82]
port 479 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[83]
port 480 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[84]
port 481 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[85]
port 482 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[86]
port 483 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[87]
port 484 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[88]
port 485 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[89]
port 486 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[8]
port 487 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[90]
port 488 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[91]
port 489 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[92]
port 490 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[93]
port 491 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[94]
port 492 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_oenb[95]
port 493 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[96]
port 494 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[97]
port 495 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_oenb[98]
port 496 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[99]
port 497 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[9]
port 498 nsew signal input
rlabel metal3 s 166334 42304 167134 42424 6 user_clock2
port 499 nsew signal input
rlabel metal3 s 166334 126896 167134 127016 6 user_irq[0]
port 500 nsew signal output
rlabel metal2 s 164882 168478 164938 169278 6 user_irq[1]
port 501 nsew signal output
rlabel metal2 s 166354 168478 166410 169278 6 user_irq[2]
port 502 nsew signal output
rlabel metal4 s 4208 2128 4528 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 34928 2128 35248 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 65648 2128 65968 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 96368 2128 96688 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 127088 2128 127408 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 157808 2128 158128 167056 6 vccd1
port 503 nsew power input
rlabel metal4 s 19568 2128 19888 167056 6 vssd1
port 504 nsew ground input
rlabel metal4 s 50288 2128 50608 167056 6 vssd1
port 504 nsew ground input
rlabel metal4 s 81008 2128 81328 167056 6 vssd1
port 504 nsew ground input
rlabel metal4 s 111728 2128 112048 167056 6 vssd1
port 504 nsew ground input
rlabel metal4 s 142448 2128 142768 167056 6 vssd1
port 504 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_ack_o
port 505 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wb_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wb_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wb_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wb_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wb_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wb_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wb_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wb_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wb_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wb_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wb_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wb_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wb_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wb_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wb_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wb_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wb_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wb_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wb_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wb_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wb_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wb_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wb_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wb_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wb_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wb_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wb_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wb_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wb_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 538 nsew signal input
rlabel metal2 s 754 0 810 800 6 wb_cyc_i
port 539 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wb_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wb_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wb_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wb_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wb_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wb_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wb_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wb_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wb_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wb_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wb_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wb_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wb_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wb_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wb_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wb_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wb_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wb_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wb_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wb_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wb_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wb_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wb_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wb_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wb_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wb_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wb_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wb_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wb_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wb_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wb_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wb_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wb_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wb_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wb_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wb_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wb_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wb_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wb_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wb_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wb_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wb_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wb_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wb_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wb_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wb_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 wb_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wb_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wb_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wb_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wb_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wb_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wb_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wb_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wb_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wb_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wb_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wb_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wb_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wb_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wb_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 604 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wb_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wb_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wb_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wb_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_stb_i
port 609 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_we_i
port 610 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 167134 169278
string LEFview TRUE
string GDS_FILE /project/openlane/sudoku_accelerator_wrapper/runs/sudoku_accelerator_wrapper/results/magic/sudoku_accelerator_wrapper.gds
string GDS_END 104759192
string GDS_START 1229370
<< end >>

