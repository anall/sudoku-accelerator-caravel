magic
tech sky130A
magscale 1 2
timestamp 1636336903
<< obsli1 >>
rect 1104 1445 180567 180625
<< obsm1 >>
rect 750 484 180579 180656
<< metal2 >>
rect 30102 182140 30158 182940
rect 90362 182140 90418 182940
rect 150622 182140 150678 182940
rect 754 0 810 800
rect 2318 0 2374 800
rect 3974 0 4030 800
rect 5630 0 5686 800
rect 7286 0 7342 800
rect 8942 0 8998 800
rect 10598 0 10654 800
rect 12254 0 12310 800
rect 13818 0 13874 800
rect 15474 0 15530 800
rect 17130 0 17186 800
rect 18786 0 18842 800
rect 20442 0 20498 800
rect 22098 0 22154 800
rect 23754 0 23810 800
rect 25318 0 25374 800
rect 26974 0 27030 800
rect 28630 0 28686 800
rect 30286 0 30342 800
rect 31942 0 31998 800
rect 33598 0 33654 800
rect 35254 0 35310 800
rect 36910 0 36966 800
rect 38474 0 38530 800
rect 40130 0 40186 800
rect 41786 0 41842 800
rect 43442 0 43498 800
rect 45098 0 45154 800
rect 46754 0 46810 800
rect 48410 0 48466 800
rect 49974 0 50030 800
rect 51630 0 51686 800
rect 53286 0 53342 800
rect 54942 0 54998 800
rect 56598 0 56654 800
rect 58254 0 58310 800
rect 59910 0 59966 800
rect 61474 0 61530 800
rect 63130 0 63186 800
rect 64786 0 64842 800
rect 66442 0 66498 800
rect 68098 0 68154 800
rect 69754 0 69810 800
rect 71410 0 71466 800
rect 73066 0 73122 800
rect 74630 0 74686 800
rect 76286 0 76342 800
rect 77942 0 77998 800
rect 79598 0 79654 800
rect 81254 0 81310 800
rect 82910 0 82966 800
rect 84566 0 84622 800
rect 86130 0 86186 800
rect 87786 0 87842 800
rect 89442 0 89498 800
rect 91098 0 91154 800
rect 92754 0 92810 800
rect 94410 0 94466 800
rect 96066 0 96122 800
rect 97630 0 97686 800
rect 99286 0 99342 800
rect 100942 0 100998 800
rect 102598 0 102654 800
rect 104254 0 104310 800
rect 105910 0 105966 800
rect 107566 0 107622 800
rect 109222 0 109278 800
rect 110786 0 110842 800
rect 112442 0 112498 800
rect 114098 0 114154 800
rect 115754 0 115810 800
rect 117410 0 117466 800
rect 119066 0 119122 800
rect 120722 0 120778 800
rect 122286 0 122342 800
rect 123942 0 123998 800
rect 125598 0 125654 800
rect 127254 0 127310 800
rect 128910 0 128966 800
rect 130566 0 130622 800
rect 132222 0 132278 800
rect 133786 0 133842 800
rect 135442 0 135498 800
rect 137098 0 137154 800
rect 138754 0 138810 800
rect 140410 0 140466 800
rect 142066 0 142122 800
rect 143722 0 143778 800
rect 145378 0 145434 800
rect 146942 0 146998 800
rect 148598 0 148654 800
rect 150254 0 150310 800
rect 151910 0 151966 800
rect 153566 0 153622 800
rect 155222 0 155278 800
rect 156878 0 156934 800
rect 158442 0 158498 800
rect 160098 0 160154 800
rect 161754 0 161810 800
rect 163410 0 163466 800
rect 165066 0 165122 800
rect 166722 0 166778 800
rect 168378 0 168434 800
rect 169942 0 169998 800
rect 171598 0 171654 800
rect 173254 0 173310 800
rect 174910 0 174966 800
rect 176566 0 176622 800
rect 178222 0 178278 800
rect 179878 0 179934 800
<< obsm2 >>
rect 756 182084 30046 182140
rect 30214 182084 90306 182140
rect 90474 182084 150566 182140
rect 150734 182084 180302 182140
rect 756 856 180302 182084
rect 866 478 2262 856
rect 2430 478 3918 856
rect 4086 478 5574 856
rect 5742 478 7230 856
rect 7398 478 8886 856
rect 9054 478 10542 856
rect 10710 478 12198 856
rect 12366 478 13762 856
rect 13930 478 15418 856
rect 15586 478 17074 856
rect 17242 478 18730 856
rect 18898 478 20386 856
rect 20554 478 22042 856
rect 22210 478 23698 856
rect 23866 478 25262 856
rect 25430 478 26918 856
rect 27086 478 28574 856
rect 28742 478 30230 856
rect 30398 478 31886 856
rect 32054 478 33542 856
rect 33710 478 35198 856
rect 35366 478 36854 856
rect 37022 478 38418 856
rect 38586 478 40074 856
rect 40242 478 41730 856
rect 41898 478 43386 856
rect 43554 478 45042 856
rect 45210 478 46698 856
rect 46866 478 48354 856
rect 48522 478 49918 856
rect 50086 478 51574 856
rect 51742 478 53230 856
rect 53398 478 54886 856
rect 55054 478 56542 856
rect 56710 478 58198 856
rect 58366 478 59854 856
rect 60022 478 61418 856
rect 61586 478 63074 856
rect 63242 478 64730 856
rect 64898 478 66386 856
rect 66554 478 68042 856
rect 68210 478 69698 856
rect 69866 478 71354 856
rect 71522 478 73010 856
rect 73178 478 74574 856
rect 74742 478 76230 856
rect 76398 478 77886 856
rect 78054 478 79542 856
rect 79710 478 81198 856
rect 81366 478 82854 856
rect 83022 478 84510 856
rect 84678 478 86074 856
rect 86242 478 87730 856
rect 87898 478 89386 856
rect 89554 478 91042 856
rect 91210 478 92698 856
rect 92866 478 94354 856
rect 94522 478 96010 856
rect 96178 478 97574 856
rect 97742 478 99230 856
rect 99398 478 100886 856
rect 101054 478 102542 856
rect 102710 478 104198 856
rect 104366 478 105854 856
rect 106022 478 107510 856
rect 107678 478 109166 856
rect 109334 478 110730 856
rect 110898 478 112386 856
rect 112554 478 114042 856
rect 114210 478 115698 856
rect 115866 478 117354 856
rect 117522 478 119010 856
rect 119178 478 120666 856
rect 120834 478 122230 856
rect 122398 478 123886 856
rect 124054 478 125542 856
rect 125710 478 127198 856
rect 127366 478 128854 856
rect 129022 478 130510 856
rect 130678 478 132166 856
rect 132334 478 133730 856
rect 133898 478 135386 856
rect 135554 478 137042 856
rect 137210 478 138698 856
rect 138866 478 140354 856
rect 140522 478 142010 856
rect 142178 478 143666 856
rect 143834 478 145322 856
rect 145490 478 146886 856
rect 147054 478 148542 856
rect 148710 478 150198 856
rect 150366 478 151854 856
rect 152022 478 153510 856
rect 153678 478 155166 856
rect 155334 478 156822 856
rect 156990 478 158386 856
rect 158554 478 160042 856
rect 160210 478 161698 856
rect 161866 478 163354 856
rect 163522 478 165010 856
rect 165178 478 166666 856
rect 166834 478 168322 856
rect 168490 478 169886 856
rect 170054 478 171542 856
rect 171710 478 173198 856
rect 173366 478 174854 856
rect 175022 478 176510 856
rect 176678 478 178166 856
rect 178334 478 179822 856
rect 179990 478 180302 856
<< obsm3 >>
rect 1117 2143 180307 180641
<< metal4 >>
rect 4208 2128 4528 180656
rect 19568 2128 19888 180656
rect 34928 2128 35248 180656
rect 50288 2128 50608 180656
rect 65648 2128 65968 180656
rect 81008 2128 81328 180656
rect 96368 2128 96688 180656
rect 111728 2128 112048 180656
rect 127088 2128 127408 180656
rect 142448 2128 142768 180656
rect 157808 2128 158128 180656
rect 173168 2128 173488 180656
<< obsm4 >>
rect 4659 4795 19488 155821
rect 19968 4795 34848 155821
rect 35328 4795 50208 155821
rect 50688 4795 65568 155821
rect 66048 4795 80928 155821
rect 81408 4795 96288 155821
rect 96768 4795 111648 155821
rect 112128 4795 127008 155821
rect 127488 4795 142368 155821
rect 142848 4795 157728 155821
rect 158208 4795 173088 155821
rect 173568 4795 174189 155821
<< labels >>
rlabel metal2 s 174910 0 174966 800 6 la_rst
port 1 nsew signal input
rlabel metal2 s 30102 182140 30158 182940 6 ser_rx
port 2 nsew signal input
rlabel metal2 s 90362 182140 90418 182940 6 ser_tx
port 3 nsew signal output
rlabel metal2 s 150622 182140 150678 182940 6 ser_tx_oeb
port 4 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 user_irq[0]
port 5 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 user_irq[1]
port 6 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 user_irq[2]
port 7 nsew signal output
rlabel metal4 s 4208 2128 4528 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 34928 2128 35248 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 65648 2128 65968 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 96368 2128 96688 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 127088 2128 127408 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 157808 2128 158128 180656 6 vccd1
port 8 nsew power input
rlabel metal4 s 19568 2128 19888 180656 6 vssd1
port 9 nsew ground input
rlabel metal4 s 50288 2128 50608 180656 6 vssd1
port 9 nsew ground input
rlabel metal4 s 81008 2128 81328 180656 6 vssd1
port 9 nsew ground input
rlabel metal4 s 111728 2128 112048 180656 6 vssd1
port 9 nsew ground input
rlabel metal4 s 142448 2128 142768 180656 6 vssd1
port 9 nsew ground input
rlabel metal4 s 173168 2128 173488 180656 6 vssd1
port 9 nsew ground input
rlabel metal2 s 754 0 810 800 6 wb_ack_o
port 10 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wb_adr_i[0]
port 11 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wb_adr_i[10]
port 12 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 wb_adr_i[11]
port 13 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 wb_adr_i[12]
port 14 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wb_adr_i[13]
port 15 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 wb_adr_i[14]
port 16 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 wb_adr_i[15]
port 17 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 wb_adr_i[16]
port 18 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 wb_adr_i[17]
port 19 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wb_adr_i[18]
port 20 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 wb_adr_i[19]
port 21 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wb_adr_i[1]
port 22 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 wb_adr_i[20]
port 23 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 wb_adr_i[21]
port 24 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 wb_adr_i[22]
port 25 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 wb_adr_i[23]
port 26 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 wb_adr_i[24]
port 27 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 wb_adr_i[25]
port 28 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 wb_adr_i[26]
port 29 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 wb_adr_i[27]
port 30 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 wb_adr_i[28]
port 31 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 wb_adr_i[29]
port 32 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wb_adr_i[2]
port 33 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 wb_adr_i[30]
port 34 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 wb_adr_i[31]
port 35 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wb_adr_i[3]
port 36 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wb_adr_i[4]
port 37 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wb_adr_i[5]
port 38 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wb_adr_i[6]
port 39 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wb_adr_i[7]
port 40 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 wb_adr_i[8]
port 41 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wb_adr_i[9]
port 42 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wb_clk_i
port 43 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wb_cyc_i
port 44 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_dat_i[0]
port 45 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wb_dat_i[10]
port 46 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wb_dat_i[11]
port 47 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 wb_dat_i[12]
port 48 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 wb_dat_i[13]
port 49 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 wb_dat_i[14]
port 50 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 wb_dat_i[15]
port 51 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wb_dat_i[16]
port 52 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 wb_dat_i[17]
port 53 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 wb_dat_i[18]
port 54 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 wb_dat_i[19]
port 55 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wb_dat_i[1]
port 56 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 wb_dat_i[20]
port 57 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 wb_dat_i[21]
port 58 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 wb_dat_i[22]
port 59 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 wb_dat_i[23]
port 60 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 wb_dat_i[24]
port 61 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 wb_dat_i[25]
port 62 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 wb_dat_i[26]
port 63 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 wb_dat_i[27]
port 64 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 wb_dat_i[28]
port 65 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 wb_dat_i[29]
port 66 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wb_dat_i[2]
port 67 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 wb_dat_i[30]
port 68 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 wb_dat_i[31]
port 69 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wb_dat_i[3]
port 70 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wb_dat_i[4]
port 71 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wb_dat_i[5]
port 72 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wb_dat_i[6]
port 73 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wb_dat_i[7]
port 74 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 wb_dat_i[8]
port 75 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wb_dat_i[9]
port 76 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wb_dat_o[0]
port 77 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 wb_dat_o[10]
port 78 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 wb_dat_o[11]
port 79 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wb_dat_o[12]
port 80 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 wb_dat_o[13]
port 81 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wb_dat_o[14]
port 82 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 wb_dat_o[15]
port 83 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 wb_dat_o[16]
port 84 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 wb_dat_o[17]
port 85 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 wb_dat_o[18]
port 86 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 wb_dat_o[19]
port 87 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 wb_dat_o[1]
port 88 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 wb_dat_o[20]
port 89 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 wb_dat_o[21]
port 90 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 wb_dat_o[22]
port 91 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 wb_dat_o[23]
port 92 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 wb_dat_o[24]
port 93 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 wb_dat_o[25]
port 94 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 wb_dat_o[26]
port 95 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 wb_dat_o[27]
port 96 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 wb_dat_o[28]
port 97 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 wb_dat_o[29]
port 98 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wb_dat_o[2]
port 99 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 wb_dat_o[30]
port 100 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 wb_dat_o[31]
port 101 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wb_dat_o[3]
port 102 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 wb_dat_o[4]
port 103 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wb_dat_o[5]
port 104 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wb_dat_o[6]
port 105 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wb_dat_o[7]
port 106 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 wb_dat_o[8]
port 107 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 wb_dat_o[9]
port 108 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wb_rst_i
port 109 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wb_sel_i[0]
port 110 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wb_sel_i[1]
port 111 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wb_sel_i[2]
port 112 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wb_sel_i[3]
port 113 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_stb_i
port 114 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb_we_i
port 115 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180796 182940
string LEFview TRUE
string GDS_FILE /project/openlane/sudoku_accelerator_wrapper/runs/sudoku_accelerator_wrapper/results/magic/sudoku_accelerator_wrapper.gds
string GDS_END 109099414
string GDS_START 1066270
<< end >>

