VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sudoku_accelerator_wrapper
  CLASS BLOCK ;
  FOREIGN sudoku_accelerator_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1315.435 BY 1326.155 ;
  PIN la_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 4.000 ;
    END
  END la_rst
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1322.155 219.330 1326.155 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 1322.155 657.710 1326.155 ;
    END
  END ser_tx
  PIN ser_tx_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 1322.155 1096.090 1326.155 ;
    END
  END ser_tx_oeb
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.790 0.000 1286.070 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1314.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1314.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1314.000 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 4.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 0.000 1022.950 4.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 4.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 0.000 819.630 4.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 0.000 1034.910 4.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 4.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 0.000 1250.190 4.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 0.000 903.350 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 0.000 1010.990 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.470 0.000 1082.750 4.000 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 0.000 1118.630 4.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 0.000 1154.510 4.000 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.990 0.000 1226.270 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.870 0.000 1262.150 4.000 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 1312.345 1309.810 1313.950 ;
        RECT 5.330 1306.905 1309.810 1309.735 ;
        RECT 5.330 1301.465 1309.810 1304.295 ;
        RECT 5.330 1296.025 1309.810 1298.855 ;
        RECT 5.330 1290.585 1309.810 1293.415 ;
        RECT 5.330 1285.145 1309.810 1287.975 ;
        RECT 5.330 1279.705 1309.810 1282.535 ;
        RECT 5.330 1274.265 1309.810 1277.095 ;
        RECT 5.330 1268.825 1309.810 1271.655 ;
        RECT 5.330 1263.385 1309.810 1266.215 ;
        RECT 5.330 1257.945 1309.810 1260.775 ;
        RECT 5.330 1252.505 1309.810 1255.335 ;
        RECT 5.330 1247.065 1309.810 1249.895 ;
        RECT 5.330 1241.625 1309.810 1244.455 ;
        RECT 5.330 1236.185 1309.810 1239.015 ;
        RECT 5.330 1230.745 1309.810 1233.575 ;
        RECT 5.330 1225.305 1309.810 1228.135 ;
        RECT 5.330 1219.865 1309.810 1222.695 ;
        RECT 5.330 1214.425 1309.810 1217.255 ;
        RECT 5.330 1208.985 1309.810 1211.815 ;
        RECT 5.330 1203.545 1309.810 1206.375 ;
        RECT 5.330 1198.105 1309.810 1200.935 ;
        RECT 5.330 1192.665 1309.810 1195.495 ;
        RECT 5.330 1187.225 1309.810 1190.055 ;
        RECT 5.330 1181.785 1309.810 1184.615 ;
        RECT 5.330 1176.345 1309.810 1179.175 ;
        RECT 5.330 1170.905 1309.810 1173.735 ;
        RECT 5.330 1165.465 1309.810 1168.295 ;
        RECT 5.330 1160.025 1309.810 1162.855 ;
        RECT 5.330 1154.585 1309.810 1157.415 ;
        RECT 5.330 1149.145 1309.810 1151.975 ;
        RECT 5.330 1143.705 1309.810 1146.535 ;
        RECT 5.330 1138.265 1309.810 1141.095 ;
        RECT 5.330 1132.825 1309.810 1135.655 ;
        RECT 5.330 1127.385 1309.810 1130.215 ;
        RECT 5.330 1121.945 1309.810 1124.775 ;
        RECT 5.330 1116.505 1309.810 1119.335 ;
        RECT 5.330 1111.065 1309.810 1113.895 ;
        RECT 5.330 1105.625 1309.810 1108.455 ;
        RECT 5.330 1100.185 1309.810 1103.015 ;
        RECT 5.330 1094.745 1309.810 1097.575 ;
        RECT 5.330 1089.305 1309.810 1092.135 ;
        RECT 5.330 1083.865 1309.810 1086.695 ;
        RECT 5.330 1078.425 1309.810 1081.255 ;
        RECT 5.330 1072.985 1309.810 1075.815 ;
        RECT 5.330 1067.545 1309.810 1070.375 ;
        RECT 5.330 1062.105 1309.810 1064.935 ;
        RECT 5.330 1056.665 1309.810 1059.495 ;
        RECT 5.330 1051.225 1309.810 1054.055 ;
        RECT 5.330 1045.785 1309.810 1048.615 ;
        RECT 5.330 1040.345 1309.810 1043.175 ;
        RECT 5.330 1034.905 1309.810 1037.735 ;
        RECT 5.330 1029.465 1309.810 1032.295 ;
        RECT 5.330 1024.025 1309.810 1026.855 ;
        RECT 5.330 1018.585 1309.810 1021.415 ;
        RECT 5.330 1013.145 1309.810 1015.975 ;
        RECT 5.330 1007.705 1309.810 1010.535 ;
        RECT 5.330 1002.265 1309.810 1005.095 ;
        RECT 5.330 996.825 1309.810 999.655 ;
        RECT 5.330 991.385 1309.810 994.215 ;
        RECT 5.330 985.945 1309.810 988.775 ;
        RECT 5.330 980.505 1309.810 983.335 ;
        RECT 5.330 975.065 1309.810 977.895 ;
        RECT 5.330 969.625 1309.810 972.455 ;
        RECT 5.330 964.185 1309.810 967.015 ;
        RECT 5.330 958.745 1309.810 961.575 ;
        RECT 5.330 953.305 1309.810 956.135 ;
        RECT 5.330 947.865 1309.810 950.695 ;
        RECT 5.330 942.425 1309.810 945.255 ;
        RECT 5.330 936.985 1309.810 939.815 ;
        RECT 5.330 931.545 1309.810 934.375 ;
        RECT 5.330 926.105 1309.810 928.935 ;
        RECT 5.330 920.665 1309.810 923.495 ;
        RECT 5.330 915.225 1309.810 918.055 ;
        RECT 5.330 909.785 1309.810 912.615 ;
        RECT 5.330 904.345 1309.810 907.175 ;
        RECT 5.330 898.905 1309.810 901.735 ;
        RECT 5.330 893.465 1309.810 896.295 ;
        RECT 5.330 888.025 1309.810 890.855 ;
        RECT 5.330 882.585 1309.810 885.415 ;
        RECT 5.330 877.145 1309.810 879.975 ;
        RECT 5.330 871.705 1309.810 874.535 ;
        RECT 5.330 866.265 1309.810 869.095 ;
        RECT 5.330 860.825 1309.810 863.655 ;
        RECT 5.330 855.385 1309.810 858.215 ;
        RECT 5.330 849.945 1309.810 852.775 ;
        RECT 5.330 844.505 1309.810 847.335 ;
        RECT 5.330 839.065 1309.810 841.895 ;
        RECT 5.330 833.625 1309.810 836.455 ;
        RECT 5.330 828.185 1309.810 831.015 ;
        RECT 5.330 822.745 1309.810 825.575 ;
        RECT 5.330 817.305 1309.810 820.135 ;
        RECT 5.330 811.865 1309.810 814.695 ;
        RECT 5.330 806.425 1309.810 809.255 ;
        RECT 5.330 800.985 1309.810 803.815 ;
        RECT 5.330 795.545 1309.810 798.375 ;
        RECT 5.330 790.105 1309.810 792.935 ;
        RECT 5.330 784.665 1309.810 787.495 ;
        RECT 5.330 779.225 1309.810 782.055 ;
        RECT 5.330 773.785 1309.810 776.615 ;
        RECT 5.330 768.345 1309.810 771.175 ;
        RECT 5.330 762.905 1309.810 765.735 ;
        RECT 5.330 757.465 1309.810 760.295 ;
        RECT 5.330 752.025 1309.810 754.855 ;
        RECT 5.330 746.585 1309.810 749.415 ;
        RECT 5.330 741.145 1309.810 743.975 ;
        RECT 5.330 735.705 1309.810 738.535 ;
        RECT 5.330 730.265 1309.810 733.095 ;
        RECT 5.330 724.825 1309.810 727.655 ;
        RECT 5.330 719.385 1309.810 722.215 ;
        RECT 5.330 713.945 1309.810 716.775 ;
        RECT 5.330 708.505 1309.810 711.335 ;
        RECT 5.330 703.065 1309.810 705.895 ;
        RECT 5.330 697.625 1309.810 700.455 ;
        RECT 5.330 692.185 1309.810 695.015 ;
        RECT 5.330 686.745 1309.810 689.575 ;
        RECT 5.330 681.305 1309.810 684.135 ;
        RECT 5.330 675.865 1309.810 678.695 ;
        RECT 5.330 670.425 1309.810 673.255 ;
        RECT 5.330 664.985 1309.810 667.815 ;
        RECT 5.330 659.545 1309.810 662.375 ;
        RECT 5.330 654.105 1309.810 656.935 ;
        RECT 5.330 648.665 1309.810 651.495 ;
        RECT 5.330 643.225 1309.810 646.055 ;
        RECT 5.330 637.785 1309.810 640.615 ;
        RECT 5.330 632.345 1309.810 635.175 ;
        RECT 5.330 626.905 1309.810 629.735 ;
        RECT 5.330 621.465 1309.810 624.295 ;
        RECT 5.330 616.025 1309.810 618.855 ;
        RECT 5.330 610.585 1309.810 613.415 ;
        RECT 5.330 605.145 1309.810 607.975 ;
        RECT 5.330 599.705 1309.810 602.535 ;
        RECT 5.330 594.265 1309.810 597.095 ;
        RECT 5.330 588.825 1309.810 591.655 ;
        RECT 5.330 583.385 1309.810 586.215 ;
        RECT 5.330 577.945 1309.810 580.775 ;
        RECT 5.330 572.505 1309.810 575.335 ;
        RECT 5.330 567.065 1309.810 569.895 ;
        RECT 5.330 561.625 1309.810 564.455 ;
        RECT 5.330 556.185 1309.810 559.015 ;
        RECT 5.330 550.745 1309.810 553.575 ;
        RECT 5.330 545.305 1309.810 548.135 ;
        RECT 5.330 539.865 1309.810 542.695 ;
        RECT 5.330 534.425 1309.810 537.255 ;
        RECT 5.330 528.985 1309.810 531.815 ;
        RECT 5.330 523.545 1309.810 526.375 ;
        RECT 5.330 518.105 1309.810 520.935 ;
        RECT 5.330 512.665 1309.810 515.495 ;
        RECT 5.330 507.225 1309.810 510.055 ;
        RECT 5.330 501.785 1309.810 504.615 ;
        RECT 5.330 496.345 1309.810 499.175 ;
        RECT 5.330 490.905 1309.810 493.735 ;
        RECT 5.330 485.465 1309.810 488.295 ;
        RECT 5.330 480.025 1309.810 482.855 ;
        RECT 5.330 474.585 1309.810 477.415 ;
        RECT 5.330 469.145 1309.810 471.975 ;
        RECT 5.330 463.705 1309.810 466.535 ;
        RECT 5.330 458.265 1309.810 461.095 ;
        RECT 5.330 452.825 1309.810 455.655 ;
        RECT 5.330 447.385 1309.810 450.215 ;
        RECT 5.330 441.945 1309.810 444.775 ;
        RECT 5.330 436.505 1309.810 439.335 ;
        RECT 5.330 431.065 1309.810 433.895 ;
        RECT 5.330 425.625 1309.810 428.455 ;
        RECT 5.330 420.185 1309.810 423.015 ;
        RECT 5.330 414.745 1309.810 417.575 ;
        RECT 5.330 409.305 1309.810 412.135 ;
        RECT 5.330 403.865 1309.810 406.695 ;
        RECT 5.330 398.425 1309.810 401.255 ;
        RECT 5.330 392.985 1309.810 395.815 ;
        RECT 5.330 387.545 1309.810 390.375 ;
        RECT 5.330 382.105 1309.810 384.935 ;
        RECT 5.330 376.665 1309.810 379.495 ;
        RECT 5.330 371.225 1309.810 374.055 ;
        RECT 5.330 365.785 1309.810 368.615 ;
        RECT 5.330 360.345 1309.810 363.175 ;
        RECT 5.330 354.905 1309.810 357.735 ;
        RECT 5.330 349.465 1309.810 352.295 ;
        RECT 5.330 344.025 1309.810 346.855 ;
        RECT 5.330 338.585 1309.810 341.415 ;
        RECT 5.330 333.145 1309.810 335.975 ;
        RECT 5.330 327.705 1309.810 330.535 ;
        RECT 5.330 322.265 1309.810 325.095 ;
        RECT 5.330 316.825 1309.810 319.655 ;
        RECT 5.330 311.385 1309.810 314.215 ;
        RECT 5.330 305.945 1309.810 308.775 ;
        RECT 5.330 300.505 1309.810 303.335 ;
        RECT 5.330 295.065 1309.810 297.895 ;
        RECT 5.330 289.625 1309.810 292.455 ;
        RECT 5.330 284.185 1309.810 287.015 ;
        RECT 5.330 278.745 1309.810 281.575 ;
        RECT 5.330 273.305 1309.810 276.135 ;
        RECT 5.330 267.865 1309.810 270.695 ;
        RECT 5.330 262.425 1309.810 265.255 ;
        RECT 5.330 256.985 1309.810 259.815 ;
        RECT 5.330 251.545 1309.810 254.375 ;
        RECT 5.330 246.105 1309.810 248.935 ;
        RECT 5.330 240.665 1309.810 243.495 ;
        RECT 5.330 235.225 1309.810 238.055 ;
        RECT 5.330 229.785 1309.810 232.615 ;
        RECT 5.330 224.345 1309.810 227.175 ;
        RECT 5.330 218.905 1309.810 221.735 ;
        RECT 5.330 213.465 1309.810 216.295 ;
        RECT 5.330 208.025 1309.810 210.855 ;
        RECT 5.330 202.585 1309.810 205.415 ;
        RECT 5.330 197.145 1309.810 199.975 ;
        RECT 5.330 191.705 1309.810 194.535 ;
        RECT 5.330 186.265 1309.810 189.095 ;
        RECT 5.330 180.825 1309.810 183.655 ;
        RECT 5.330 175.385 1309.810 178.215 ;
        RECT 5.330 169.945 1309.810 172.775 ;
        RECT 5.330 164.505 1309.810 167.335 ;
        RECT 5.330 159.065 1309.810 161.895 ;
        RECT 5.330 153.625 1309.810 156.455 ;
        RECT 5.330 148.185 1309.810 151.015 ;
        RECT 5.330 142.745 1309.810 145.575 ;
        RECT 5.330 137.305 1309.810 140.135 ;
        RECT 5.330 131.865 1309.810 134.695 ;
        RECT 5.330 126.425 1309.810 129.255 ;
        RECT 5.330 120.985 1309.810 123.815 ;
        RECT 5.330 115.545 1309.810 118.375 ;
        RECT 5.330 110.105 1309.810 112.935 ;
        RECT 5.330 104.665 1309.810 107.495 ;
        RECT 5.330 99.225 1309.810 102.055 ;
        RECT 5.330 93.785 1309.810 96.615 ;
        RECT 5.330 88.345 1309.810 91.175 ;
        RECT 5.330 82.905 1309.810 85.735 ;
        RECT 5.330 77.465 1309.810 80.295 ;
        RECT 5.330 72.025 1309.810 74.855 ;
        RECT 5.330 66.585 1309.810 69.415 ;
        RECT 5.330 61.145 1309.810 63.975 ;
        RECT 5.330 55.705 1309.810 58.535 ;
        RECT 5.330 50.265 1309.810 53.095 ;
        RECT 5.330 44.825 1309.810 47.655 ;
        RECT 5.330 39.385 1309.810 42.215 ;
        RECT 5.330 33.945 1309.810 36.775 ;
        RECT 5.330 28.505 1309.810 31.335 ;
        RECT 5.330 23.065 1309.810 25.895 ;
        RECT 5.330 17.625 1309.810 20.455 ;
        RECT 5.330 12.185 1309.810 15.015 ;
      LAYER li1 ;
        RECT 5.520 6.885 1309.620 1313.845 ;
      LAYER met1 ;
        RECT 5.520 6.840 1310.010 1314.000 ;
      LAYER met2 ;
        RECT 6.080 1321.875 218.770 1322.155 ;
        RECT 219.610 1321.875 657.150 1322.155 ;
        RECT 657.990 1321.875 1095.530 1322.155 ;
        RECT 1096.370 1321.875 1309.980 1322.155 ;
        RECT 6.080 4.280 1309.980 1321.875 ;
        RECT 6.630 3.670 17.750 4.280 ;
        RECT 18.590 3.670 29.710 4.280 ;
        RECT 30.550 3.670 41.670 4.280 ;
        RECT 42.510 3.670 53.630 4.280 ;
        RECT 54.470 3.670 65.590 4.280 ;
        RECT 66.430 3.670 77.550 4.280 ;
        RECT 78.390 3.670 89.510 4.280 ;
        RECT 90.350 3.670 101.470 4.280 ;
        RECT 102.310 3.670 113.430 4.280 ;
        RECT 114.270 3.670 125.390 4.280 ;
        RECT 126.230 3.670 137.350 4.280 ;
        RECT 138.190 3.670 149.310 4.280 ;
        RECT 150.150 3.670 161.270 4.280 ;
        RECT 162.110 3.670 173.230 4.280 ;
        RECT 174.070 3.670 185.190 4.280 ;
        RECT 186.030 3.670 197.150 4.280 ;
        RECT 197.990 3.670 209.110 4.280 ;
        RECT 209.950 3.670 221.070 4.280 ;
        RECT 221.910 3.670 233.030 4.280 ;
        RECT 233.870 3.670 244.990 4.280 ;
        RECT 245.830 3.670 256.950 4.280 ;
        RECT 257.790 3.670 268.910 4.280 ;
        RECT 269.750 3.670 280.870 4.280 ;
        RECT 281.710 3.670 292.830 4.280 ;
        RECT 293.670 3.670 304.790 4.280 ;
        RECT 305.630 3.670 316.750 4.280 ;
        RECT 317.590 3.670 328.710 4.280 ;
        RECT 329.550 3.670 340.670 4.280 ;
        RECT 341.510 3.670 352.630 4.280 ;
        RECT 353.470 3.670 364.590 4.280 ;
        RECT 365.430 3.670 376.550 4.280 ;
        RECT 377.390 3.670 388.510 4.280 ;
        RECT 389.350 3.670 400.470 4.280 ;
        RECT 401.310 3.670 412.430 4.280 ;
        RECT 413.270 3.670 424.390 4.280 ;
        RECT 425.230 3.670 436.350 4.280 ;
        RECT 437.190 3.670 448.310 4.280 ;
        RECT 449.150 3.670 460.270 4.280 ;
        RECT 461.110 3.670 472.230 4.280 ;
        RECT 473.070 3.670 484.190 4.280 ;
        RECT 485.030 3.670 496.150 4.280 ;
        RECT 496.990 3.670 508.110 4.280 ;
        RECT 508.950 3.670 520.070 4.280 ;
        RECT 520.910 3.670 532.030 4.280 ;
        RECT 532.870 3.670 543.990 4.280 ;
        RECT 544.830 3.670 555.950 4.280 ;
        RECT 556.790 3.670 567.910 4.280 ;
        RECT 568.750 3.670 579.870 4.280 ;
        RECT 580.710 3.670 591.830 4.280 ;
        RECT 592.670 3.670 603.790 4.280 ;
        RECT 604.630 3.670 615.750 4.280 ;
        RECT 616.590 3.670 627.710 4.280 ;
        RECT 628.550 3.670 639.670 4.280 ;
        RECT 640.510 3.670 651.630 4.280 ;
        RECT 652.470 3.670 663.590 4.280 ;
        RECT 664.430 3.670 675.550 4.280 ;
        RECT 676.390 3.670 687.510 4.280 ;
        RECT 688.350 3.670 699.470 4.280 ;
        RECT 700.310 3.670 711.430 4.280 ;
        RECT 712.270 3.670 723.390 4.280 ;
        RECT 724.230 3.670 735.350 4.280 ;
        RECT 736.190 3.670 747.310 4.280 ;
        RECT 748.150 3.670 759.270 4.280 ;
        RECT 760.110 3.670 771.230 4.280 ;
        RECT 772.070 3.670 783.190 4.280 ;
        RECT 784.030 3.670 795.150 4.280 ;
        RECT 795.990 3.670 807.110 4.280 ;
        RECT 807.950 3.670 819.070 4.280 ;
        RECT 819.910 3.670 831.030 4.280 ;
        RECT 831.870 3.670 842.990 4.280 ;
        RECT 843.830 3.670 854.950 4.280 ;
        RECT 855.790 3.670 866.910 4.280 ;
        RECT 867.750 3.670 878.870 4.280 ;
        RECT 879.710 3.670 890.830 4.280 ;
        RECT 891.670 3.670 902.790 4.280 ;
        RECT 903.630 3.670 914.750 4.280 ;
        RECT 915.590 3.670 926.710 4.280 ;
        RECT 927.550 3.670 938.670 4.280 ;
        RECT 939.510 3.670 950.630 4.280 ;
        RECT 951.470 3.670 962.590 4.280 ;
        RECT 963.430 3.670 974.550 4.280 ;
        RECT 975.390 3.670 986.510 4.280 ;
        RECT 987.350 3.670 998.470 4.280 ;
        RECT 999.310 3.670 1010.430 4.280 ;
        RECT 1011.270 3.670 1022.390 4.280 ;
        RECT 1023.230 3.670 1034.350 4.280 ;
        RECT 1035.190 3.670 1046.310 4.280 ;
        RECT 1047.150 3.670 1058.270 4.280 ;
        RECT 1059.110 3.670 1070.230 4.280 ;
        RECT 1071.070 3.670 1082.190 4.280 ;
        RECT 1083.030 3.670 1094.150 4.280 ;
        RECT 1094.990 3.670 1106.110 4.280 ;
        RECT 1106.950 3.670 1118.070 4.280 ;
        RECT 1118.910 3.670 1130.030 4.280 ;
        RECT 1130.870 3.670 1141.990 4.280 ;
        RECT 1142.830 3.670 1153.950 4.280 ;
        RECT 1154.790 3.670 1165.910 4.280 ;
        RECT 1166.750 3.670 1177.870 4.280 ;
        RECT 1178.710 3.670 1189.830 4.280 ;
        RECT 1190.670 3.670 1201.790 4.280 ;
        RECT 1202.630 3.670 1213.750 4.280 ;
        RECT 1214.590 3.670 1225.710 4.280 ;
        RECT 1226.550 3.670 1237.670 4.280 ;
        RECT 1238.510 3.670 1249.630 4.280 ;
        RECT 1250.470 3.670 1261.590 4.280 ;
        RECT 1262.430 3.670 1273.550 4.280 ;
        RECT 1274.390 3.670 1285.510 4.280 ;
        RECT 1286.350 3.670 1297.470 4.280 ;
        RECT 1298.310 3.670 1309.430 4.280 ;
      LAYER met3 ;
        RECT 10.185 9.015 1299.895 1313.925 ;
      LAYER met4 ;
        RECT 49.055 10.240 97.440 1311.545 ;
        RECT 99.840 10.240 174.240 1311.545 ;
        RECT 176.640 10.240 251.040 1311.545 ;
        RECT 253.440 10.240 327.840 1311.545 ;
        RECT 330.240 10.240 404.640 1311.545 ;
        RECT 407.040 10.240 481.440 1311.545 ;
        RECT 483.840 10.240 558.240 1311.545 ;
        RECT 560.640 10.240 635.040 1311.545 ;
        RECT 637.440 10.240 711.840 1311.545 ;
        RECT 714.240 10.240 788.640 1311.545 ;
        RECT 791.040 10.240 865.440 1311.545 ;
        RECT 867.840 10.240 942.240 1311.545 ;
        RECT 944.640 10.240 1019.040 1311.545 ;
        RECT 1021.440 10.240 1065.985 1311.545 ;
        RECT 49.055 9.015 1065.985 10.240 ;
  END
END sudoku_accelerator_wrapper
END LIBRARY

