magic
tech sky130A
magscale 1 2
timestamp 1635789796
<< nwell >>
rect 1066 262469 261962 262790
rect 1066 261381 261962 261947
rect 1066 260293 261962 260859
rect 1066 259205 261962 259771
rect 1066 258117 261962 258683
rect 1066 257029 261962 257595
rect 1066 255941 261962 256507
rect 1066 254853 261962 255419
rect 1066 253765 261962 254331
rect 1066 252677 261962 253243
rect 1066 251589 261962 252155
rect 1066 250501 261962 251067
rect 1066 249413 261962 249979
rect 1066 248325 261962 248891
rect 1066 247237 261962 247803
rect 1066 246149 261962 246715
rect 1066 245061 261962 245627
rect 1066 243973 261962 244539
rect 1066 242885 261962 243451
rect 1066 241797 261962 242363
rect 1066 240709 261962 241275
rect 1066 239621 261962 240187
rect 1066 238533 261962 239099
rect 1066 237445 261962 238011
rect 1066 236357 261962 236923
rect 1066 235269 261962 235835
rect 1066 234181 261962 234747
rect 1066 233093 261962 233659
rect 1066 232005 261962 232571
rect 1066 230917 261962 231483
rect 1066 229829 261962 230395
rect 1066 228741 261962 229307
rect 1066 227653 261962 228219
rect 1066 226565 261962 227131
rect 1066 225477 261962 226043
rect 1066 224389 261962 224955
rect 1066 223301 261962 223867
rect 1066 222213 261962 222779
rect 1066 221125 261962 221691
rect 1066 220037 261962 220603
rect 1066 218949 261962 219515
rect 1066 217861 261962 218427
rect 1066 216773 261962 217339
rect 1066 215685 261962 216251
rect 1066 214597 261962 215163
rect 1066 213509 261962 214075
rect 1066 212421 261962 212987
rect 1066 211333 261962 211899
rect 1066 210245 261962 210811
rect 1066 209157 261962 209723
rect 1066 208069 261962 208635
rect 1066 206981 261962 207547
rect 1066 205893 261962 206459
rect 1066 204805 261962 205371
rect 1066 203717 261962 204283
rect 1066 202629 261962 203195
rect 1066 201541 261962 202107
rect 1066 200453 261962 201019
rect 1066 199365 261962 199931
rect 1066 198277 261962 198843
rect 1066 197189 261962 197755
rect 1066 196101 261962 196667
rect 1066 195013 261962 195579
rect 1066 193925 261962 194491
rect 1066 192837 261962 193403
rect 1066 191749 261962 192315
rect 1066 190661 261962 191227
rect 1066 189573 261962 190139
rect 1066 188485 261962 189051
rect 1066 187397 261962 187963
rect 1066 186309 261962 186875
rect 1066 185221 261962 185787
rect 1066 184133 261962 184699
rect 1066 183045 261962 183611
rect 1066 181957 261962 182523
rect 1066 180869 261962 181435
rect 1066 179781 261962 180347
rect 1066 178693 261962 179259
rect 1066 177605 261962 178171
rect 1066 176517 261962 177083
rect 1066 175429 261962 175995
rect 1066 174341 261962 174907
rect 1066 173253 261962 173819
rect 1066 172165 261962 172731
rect 1066 171077 261962 171643
rect 1066 169989 261962 170555
rect 1066 168901 261962 169467
rect 1066 167813 261962 168379
rect 1066 166725 261962 167291
rect 1066 165637 261962 166203
rect 1066 164549 261962 165115
rect 1066 163461 261962 164027
rect 1066 162373 261962 162939
rect 1066 161285 261962 161851
rect 1066 160197 261962 160763
rect 1066 159109 261962 159675
rect 1066 158021 261962 158587
rect 1066 156933 261962 157499
rect 1066 155845 261962 156411
rect 1066 154757 261962 155323
rect 1066 153669 261962 154235
rect 1066 152581 261962 153147
rect 1066 151493 261962 152059
rect 1066 150405 261962 150971
rect 1066 149317 261962 149883
rect 1066 148229 261962 148795
rect 1066 147141 261962 147707
rect 1066 146053 261962 146619
rect 1066 144965 261962 145531
rect 1066 143877 261962 144443
rect 1066 142789 261962 143355
rect 1066 141701 261962 142267
rect 1066 140613 261962 141179
rect 1066 139525 261962 140091
rect 1066 138437 261962 139003
rect 1066 137349 261962 137915
rect 1066 136261 261962 136827
rect 1066 135173 261962 135739
rect 1066 134085 261962 134651
rect 1066 132997 261962 133563
rect 1066 131909 261962 132475
rect 1066 130821 261962 131387
rect 1066 129733 261962 130299
rect 1066 128645 261962 129211
rect 1066 127557 261962 128123
rect 1066 126469 261962 127035
rect 1066 125381 261962 125947
rect 1066 124293 261962 124859
rect 1066 123205 261962 123771
rect 1066 122117 261962 122683
rect 1066 121029 261962 121595
rect 1066 119941 261962 120507
rect 1066 118853 261962 119419
rect 1066 117765 261962 118331
rect 1066 116677 261962 117243
rect 1066 115589 261962 116155
rect 1066 114501 261962 115067
rect 1066 113413 261962 113979
rect 1066 112325 261962 112891
rect 1066 111237 261962 111803
rect 1066 110149 261962 110715
rect 1066 109061 261962 109627
rect 1066 107973 261962 108539
rect 1066 106885 261962 107451
rect 1066 105797 261962 106363
rect 1066 104709 261962 105275
rect 1066 103621 261962 104187
rect 1066 102533 261962 103099
rect 1066 101445 261962 102011
rect 1066 100357 261962 100923
rect 1066 99269 261962 99835
rect 1066 98181 261962 98747
rect 1066 97093 261962 97659
rect 1066 96005 261962 96571
rect 1066 94917 261962 95483
rect 1066 93829 261962 94395
rect 1066 92741 261962 93307
rect 1066 91653 261962 92219
rect 1066 90565 261962 91131
rect 1066 89477 261962 90043
rect 1066 88389 261962 88955
rect 1066 87301 261962 87867
rect 1066 86213 261962 86779
rect 1066 85125 261962 85691
rect 1066 84037 261962 84603
rect 1066 82949 261962 83515
rect 1066 81861 261962 82427
rect 1066 80773 261962 81339
rect 1066 79685 261962 80251
rect 1066 78597 261962 79163
rect 1066 77509 261962 78075
rect 1066 76421 261962 76987
rect 1066 75333 261962 75899
rect 1066 74245 261962 74811
rect 1066 73157 261962 73723
rect 1066 72069 261962 72635
rect 1066 70981 261962 71547
rect 1066 69893 261962 70459
rect 1066 68805 261962 69371
rect 1066 67717 261962 68283
rect 1066 66629 261962 67195
rect 1066 65541 261962 66107
rect 1066 64453 261962 65019
rect 1066 63365 261962 63931
rect 1066 62277 261962 62843
rect 1066 61189 261962 61755
rect 1066 60101 261962 60667
rect 1066 59013 261962 59579
rect 1066 57925 261962 58491
rect 1066 56837 261962 57403
rect 1066 55749 261962 56315
rect 1066 54661 261962 55227
rect 1066 53573 261962 54139
rect 1066 52485 261962 53051
rect 1066 51397 261962 51963
rect 1066 50309 261962 50875
rect 1066 49221 261962 49787
rect 1066 48133 261962 48699
rect 1066 47045 261962 47611
rect 1066 45957 261962 46523
rect 1066 44869 261962 45435
rect 1066 43781 261962 44347
rect 1066 42693 261962 43259
rect 1066 41605 261962 42171
rect 1066 40517 261962 41083
rect 1066 39429 261962 39995
rect 1066 38341 261962 38907
rect 1066 37253 261962 37819
rect 1066 36165 261962 36731
rect 1066 35077 261962 35643
rect 1066 33989 261962 34555
rect 1066 32901 261962 33467
rect 1066 31813 261962 32379
rect 1066 30725 261962 31291
rect 1066 29637 261962 30203
rect 1066 28549 261962 29115
rect 1066 27461 261962 28027
rect 1066 26373 261962 26939
rect 1066 25285 261962 25851
rect 1066 24197 261962 24763
rect 1066 23109 261962 23675
rect 1066 22021 261962 22587
rect 1066 20933 261962 21499
rect 1066 19845 261962 20411
rect 1066 18757 261962 19323
rect 1066 17669 261962 18235
rect 1066 16581 261962 17147
rect 1066 15493 261962 16059
rect 1066 14405 261962 14971
rect 1066 13317 261962 13883
rect 1066 12229 261962 12795
rect 1066 11141 261962 11707
rect 1066 10053 261962 10619
rect 1066 8965 261962 9531
rect 1066 7877 261962 8443
rect 1066 6789 261962 7355
rect 1066 5701 261962 6267
rect 1066 4613 261962 5179
rect 1066 3525 261962 4091
rect 1066 2437 261962 3003
<< obsli1 >>
rect 1104 1377 261924 262769
<< obsm1 >>
rect 1104 1368 262002 262800
<< metal2 >>
rect 43810 264431 43866 265231
rect 131486 264431 131542 265231
rect 219162 264431 219218 265231
rect 1214 0 1270 800
rect 3606 0 3662 800
rect 5998 0 6054 800
rect 8390 0 8446 800
rect 10782 0 10838 800
rect 13174 0 13230 800
rect 15566 0 15622 800
rect 17958 0 18014 800
rect 20350 0 20406 800
rect 22742 0 22798 800
rect 25134 0 25190 800
rect 27526 0 27582 800
rect 29918 0 29974 800
rect 32310 0 32366 800
rect 34702 0 34758 800
rect 37094 0 37150 800
rect 39486 0 39542 800
rect 41878 0 41934 800
rect 44270 0 44326 800
rect 46662 0 46718 800
rect 49054 0 49110 800
rect 51446 0 51502 800
rect 53838 0 53894 800
rect 56230 0 56286 800
rect 58622 0 58678 800
rect 61014 0 61070 800
rect 63406 0 63462 800
rect 65798 0 65854 800
rect 68190 0 68246 800
rect 70582 0 70638 800
rect 72974 0 73030 800
rect 75366 0 75422 800
rect 77758 0 77814 800
rect 80150 0 80206 800
rect 82542 0 82598 800
rect 84934 0 84990 800
rect 87326 0 87382 800
rect 89718 0 89774 800
rect 92110 0 92166 800
rect 94502 0 94558 800
rect 96894 0 96950 800
rect 99286 0 99342 800
rect 101678 0 101734 800
rect 104070 0 104126 800
rect 106462 0 106518 800
rect 108854 0 108910 800
rect 111246 0 111302 800
rect 113638 0 113694 800
rect 116030 0 116086 800
rect 118422 0 118478 800
rect 120814 0 120870 800
rect 123206 0 123262 800
rect 125598 0 125654 800
rect 127990 0 128046 800
rect 130382 0 130438 800
rect 132774 0 132830 800
rect 135166 0 135222 800
rect 137558 0 137614 800
rect 139950 0 140006 800
rect 142342 0 142398 800
rect 144734 0 144790 800
rect 147126 0 147182 800
rect 149518 0 149574 800
rect 151910 0 151966 800
rect 154302 0 154358 800
rect 156694 0 156750 800
rect 159086 0 159142 800
rect 161478 0 161534 800
rect 163870 0 163926 800
rect 166262 0 166318 800
rect 168654 0 168710 800
rect 171046 0 171102 800
rect 173438 0 173494 800
rect 175830 0 175886 800
rect 178222 0 178278 800
rect 180614 0 180670 800
rect 183006 0 183062 800
rect 185398 0 185454 800
rect 187790 0 187846 800
rect 190182 0 190238 800
rect 192574 0 192630 800
rect 194966 0 195022 800
rect 197358 0 197414 800
rect 199750 0 199806 800
rect 202142 0 202198 800
rect 204534 0 204590 800
rect 206926 0 206982 800
rect 209318 0 209374 800
rect 211710 0 211766 800
rect 214102 0 214158 800
rect 216494 0 216550 800
rect 218886 0 218942 800
rect 221278 0 221334 800
rect 223670 0 223726 800
rect 226062 0 226118 800
rect 228454 0 228510 800
rect 230846 0 230902 800
rect 233238 0 233294 800
rect 235630 0 235686 800
rect 238022 0 238078 800
rect 240414 0 240470 800
rect 242806 0 242862 800
rect 245198 0 245254 800
rect 247590 0 247646 800
rect 249982 0 250038 800
rect 252374 0 252430 800
rect 254766 0 254822 800
rect 257158 0 257214 800
rect 259550 0 259606 800
rect 261942 0 261998 800
<< obsm2 >>
rect 1216 264375 43754 264431
rect 43922 264375 131430 264431
rect 131598 264375 219106 264431
rect 219274 264375 261996 264431
rect 1216 856 261996 264375
rect 1326 734 3550 856
rect 3718 734 5942 856
rect 6110 734 8334 856
rect 8502 734 10726 856
rect 10894 734 13118 856
rect 13286 734 15510 856
rect 15678 734 17902 856
rect 18070 734 20294 856
rect 20462 734 22686 856
rect 22854 734 25078 856
rect 25246 734 27470 856
rect 27638 734 29862 856
rect 30030 734 32254 856
rect 32422 734 34646 856
rect 34814 734 37038 856
rect 37206 734 39430 856
rect 39598 734 41822 856
rect 41990 734 44214 856
rect 44382 734 46606 856
rect 46774 734 48998 856
rect 49166 734 51390 856
rect 51558 734 53782 856
rect 53950 734 56174 856
rect 56342 734 58566 856
rect 58734 734 60958 856
rect 61126 734 63350 856
rect 63518 734 65742 856
rect 65910 734 68134 856
rect 68302 734 70526 856
rect 70694 734 72918 856
rect 73086 734 75310 856
rect 75478 734 77702 856
rect 77870 734 80094 856
rect 80262 734 82486 856
rect 82654 734 84878 856
rect 85046 734 87270 856
rect 87438 734 89662 856
rect 89830 734 92054 856
rect 92222 734 94446 856
rect 94614 734 96838 856
rect 97006 734 99230 856
rect 99398 734 101622 856
rect 101790 734 104014 856
rect 104182 734 106406 856
rect 106574 734 108798 856
rect 108966 734 111190 856
rect 111358 734 113582 856
rect 113750 734 115974 856
rect 116142 734 118366 856
rect 118534 734 120758 856
rect 120926 734 123150 856
rect 123318 734 125542 856
rect 125710 734 127934 856
rect 128102 734 130326 856
rect 130494 734 132718 856
rect 132886 734 135110 856
rect 135278 734 137502 856
rect 137670 734 139894 856
rect 140062 734 142286 856
rect 142454 734 144678 856
rect 144846 734 147070 856
rect 147238 734 149462 856
rect 149630 734 151854 856
rect 152022 734 154246 856
rect 154414 734 156638 856
rect 156806 734 159030 856
rect 159198 734 161422 856
rect 161590 734 163814 856
rect 163982 734 166206 856
rect 166374 734 168598 856
rect 168766 734 170990 856
rect 171158 734 173382 856
rect 173550 734 175774 856
rect 175942 734 178166 856
rect 178334 734 180558 856
rect 180726 734 182950 856
rect 183118 734 185342 856
rect 185510 734 187734 856
rect 187902 734 190126 856
rect 190294 734 192518 856
rect 192686 734 194910 856
rect 195078 734 197302 856
rect 197470 734 199694 856
rect 199862 734 202086 856
rect 202254 734 204478 856
rect 204646 734 206870 856
rect 207038 734 209262 856
rect 209430 734 211654 856
rect 211822 734 214046 856
rect 214214 734 216438 856
rect 216606 734 218830 856
rect 218998 734 221222 856
rect 221390 734 223614 856
rect 223782 734 226006 856
rect 226174 734 228398 856
rect 228566 734 230790 856
rect 230958 734 233182 856
rect 233350 734 235574 856
rect 235742 734 237966 856
rect 238134 734 240358 856
rect 240526 734 242750 856
rect 242918 734 245142 856
rect 245310 734 247534 856
rect 247702 734 249926 856
rect 250094 734 252318 856
rect 252486 734 254710 856
rect 254878 734 257102 856
rect 257270 734 259494 856
rect 259662 734 261886 856
<< obsm3 >>
rect 2037 1803 259979 262785
<< metal4 >>
rect 4208 2128 4528 262800
rect 19568 2128 19888 262800
rect 34928 2128 35248 262800
rect 50288 2128 50608 262800
rect 65648 2128 65968 262800
rect 81008 2128 81328 262800
rect 96368 2128 96688 262800
rect 111728 2128 112048 262800
rect 127088 2128 127408 262800
rect 142448 2128 142768 262800
rect 157808 2128 158128 262800
rect 173168 2128 173488 262800
rect 188528 2128 188848 262800
rect 203888 2128 204208 262800
rect 219248 2128 219568 262800
rect 234608 2128 234928 262800
rect 249968 2128 250288 262800
<< obsm4 >>
rect 9811 2048 19488 262309
rect 19968 2048 34848 262309
rect 35328 2048 50208 262309
rect 50688 2048 65568 262309
rect 66048 2048 80928 262309
rect 81408 2048 96288 262309
rect 96768 2048 111648 262309
rect 112128 2048 127008 262309
rect 127488 2048 142368 262309
rect 142848 2048 157728 262309
rect 158208 2048 173088 262309
rect 173568 2048 188448 262309
rect 188928 2048 203808 262309
rect 204288 2048 213197 262309
rect 9811 1803 213197 2048
<< labels >>
rlabel metal2 s 254766 0 254822 800 6 la_rst
port 1 nsew signal input
rlabel metal2 s 43810 264431 43866 265231 6 ser_rx
port 2 nsew signal input
rlabel metal2 s 131486 264431 131542 265231 6 ser_tx
port 3 nsew signal output
rlabel metal2 s 219162 264431 219218 265231 6 ser_tx_oeb
port 4 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 user_irq[0]
port 5 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 user_irq[1]
port 6 nsew signal output
rlabel metal2 s 261942 0 261998 800 6 user_irq[2]
port 7 nsew signal output
rlabel metal4 s 4208 2128 4528 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 34928 2128 35248 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 65648 2128 65968 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 96368 2128 96688 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 127088 2128 127408 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 157808 2128 158128 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 188528 2128 188848 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 219248 2128 219568 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 249968 2128 250288 262800 6 vccd1
port 8 nsew power input
rlabel metal4 s 19568 2128 19888 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 50288 2128 50608 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 81008 2128 81328 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 111728 2128 112048 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 142448 2128 142768 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 173168 2128 173488 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 203888 2128 204208 262800 6 vssd1
port 9 nsew ground input
rlabel metal4 s 234608 2128 234928 262800 6 vssd1
port 9 nsew ground input
rlabel metal2 s 1214 0 1270 800 6 wb_ack_o
port 10 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wb_adr_i[0]
port 11 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 wb_adr_i[10]
port 12 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 wb_adr_i[11]
port 13 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wb_adr_i[12]
port 14 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 wb_adr_i[13]
port 15 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 wb_adr_i[14]
port 16 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 wb_adr_i[15]
port 17 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 wb_adr_i[16]
port 18 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 wb_adr_i[17]
port 19 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 wb_adr_i[18]
port 20 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 wb_adr_i[19]
port 21 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wb_adr_i[1]
port 22 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 wb_adr_i[20]
port 23 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 wb_adr_i[21]
port 24 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 wb_adr_i[22]
port 25 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 wb_adr_i[23]
port 26 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 wb_adr_i[24]
port 27 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 wb_adr_i[25]
port 28 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 wb_adr_i[26]
port 29 nsew signal input
rlabel metal2 s 218886 0 218942 800 6 wb_adr_i[27]
port 30 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 wb_adr_i[28]
port 31 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 wb_adr_i[29]
port 32 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wb_adr_i[2]
port 33 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 wb_adr_i[30]
port 34 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 wb_adr_i[31]
port 35 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wb_adr_i[3]
port 36 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wb_adr_i[4]
port 37 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wb_adr_i[5]
port 38 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 wb_adr_i[6]
port 39 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 wb_adr_i[7]
port 40 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wb_adr_i[8]
port 41 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 wb_adr_i[9]
port 42 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wb_clk_i
port 43 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_cyc_i
port 44 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wb_dat_i[0]
port 45 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wb_dat_i[10]
port 46 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 wb_dat_i[11]
port 47 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 wb_dat_i[12]
port 48 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 wb_dat_i[13]
port 49 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 wb_dat_i[14]
port 50 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 wb_dat_i[15]
port 51 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 wb_dat_i[16]
port 52 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 wb_dat_i[17]
port 53 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 wb_dat_i[18]
port 54 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 wb_dat_i[19]
port 55 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wb_dat_i[1]
port 56 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 wb_dat_i[20]
port 57 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 wb_dat_i[21]
port 58 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 wb_dat_i[22]
port 59 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 wb_dat_i[23]
port 60 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 wb_dat_i[24]
port 61 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 wb_dat_i[25]
port 62 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 wb_dat_i[26]
port 63 nsew signal input
rlabel metal2 s 221278 0 221334 800 6 wb_dat_i[27]
port 64 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 wb_dat_i[28]
port 65 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 wb_dat_i[29]
port 66 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wb_dat_i[2]
port 67 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 wb_dat_i[30]
port 68 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 wb_dat_i[31]
port 69 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wb_dat_i[3]
port 70 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wb_dat_i[4]
port 71 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wb_dat_i[5]
port 72 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wb_dat_i[6]
port 73 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wb_dat_i[7]
port 74 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wb_dat_i[8]
port 75 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 wb_dat_i[9]
port 76 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wb_dat_o[0]
port 77 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 wb_dat_o[10]
port 78 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 wb_dat_o[11]
port 79 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wb_dat_o[12]
port 80 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 wb_dat_o[13]
port 81 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 wb_dat_o[14]
port 82 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 wb_dat_o[15]
port 83 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 wb_dat_o[16]
port 84 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 wb_dat_o[17]
port 85 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 wb_dat_o[18]
port 86 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 wb_dat_o[19]
port 87 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 wb_dat_o[1]
port 88 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 wb_dat_o[20]
port 89 nsew signal output
rlabel metal2 s 180614 0 180670 800 6 wb_dat_o[21]
port 90 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 wb_dat_o[22]
port 91 nsew signal output
rlabel metal2 s 194966 0 195022 800 6 wb_dat_o[23]
port 92 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 wb_dat_o[24]
port 93 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 wb_dat_o[25]
port 94 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 wb_dat_o[26]
port 95 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 wb_dat_o[27]
port 96 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 wb_dat_o[28]
port 97 nsew signal output
rlabel metal2 s 238022 0 238078 800 6 wb_dat_o[29]
port 98 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 wb_dat_o[2]
port 99 nsew signal output
rlabel metal2 s 245198 0 245254 800 6 wb_dat_o[30]
port 100 nsew signal output
rlabel metal2 s 252374 0 252430 800 6 wb_dat_o[31]
port 101 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 wb_dat_o[3]
port 102 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wb_dat_o[4]
port 103 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 wb_dat_o[5]
port 104 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 wb_dat_o[6]
port 105 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 wb_dat_o[7]
port 106 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 wb_dat_o[8]
port 107 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 wb_dat_o[9]
port 108 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wb_rst_i
port 109 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wb_sel_i[0]
port 110 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wb_sel_i[1]
port 111 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wb_sel_i[2]
port 112 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wb_sel_i[3]
port 113 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wb_stb_i
port 114 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_we_i
port 115 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 263087 265231
string LEFview TRUE
string GDS_FILE /project/openlane/sudoku_accelerator_wrapper/runs/sudoku_accelerator_wrapper/results/magic/sudoku_accelerator_wrapper.gds
string GDS_END 124935646
string GDS_START 1393548
<< end >>

